library verilog;
use verilog.vl_types.all;
entity IF_tb is
end IF_tb;
