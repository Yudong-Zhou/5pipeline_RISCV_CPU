//******************************************************************************
// Author:Zhou Yudong
// ALU.v
//******************************************************************************
module ALU (
	// Outputs
	ALUResult,
	// Inputs
	ALUCode, A, B);
	input [3:0]	ALUCode;				// Operation select
	input [31:0]	A, B;
	output [31:0]	ALUResult;
	
// Decoded ALU operation select (ALUsel) signals
  parameter	 alu_add=  4'b0000;
  parameter	 alu_sub=  4'b0001;
  parameter	 alu_lui=  4'b0010;
  parameter	 alu_and=  4'b0011;
  parameter	 alu_xor=  4'b0100;
  parameter	 alu_or =  4'b0101;
  parameter 	alu_sll=  4'b0110;
  parameter	 alu_srl=  4'b0111;
  parameter	 alu_sra=  4'b1000;
  parameter	 alu_slt=  4'b1001;
  parameter	 alu_sltu= 4'b1010; 	

  wire Binvert;
  reg Binvert_32bits;
  assign Binvert = ~(ALUCode == 0);
  always@(*) begin
    if(~Binvert) Binvert_32bits = {31'b0,Binvert};
    else Binvert_32bits = {31'b1,Binvert};
  end
  
  
  
  
  
endmodule