library verilog;
use verilog.vl_types.all;
entity Decode_tb is
end Decode_tb;
